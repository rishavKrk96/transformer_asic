##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Sun Mar 19 01:54:55 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 766.400000 BY 765.200000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 357.300000 0.600000 357.500000 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 357.700000 0.600000 357.900000 ;
    END
  END clk2
  PIN mem_in1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 393.700000 0.600000 393.900000 ;
    END
  END mem_in1[31]
  PIN mem_in1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 393.300000 0.600000 393.500000 ;
    END
  END mem_in1[30]
  PIN mem_in1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.900000 0.600000 393.100000 ;
    END
  END mem_in1[29]
  PIN mem_in1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.500000 0.600000 392.700000 ;
    END
  END mem_in1[28]
  PIN mem_in1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.100000 0.600000 392.300000 ;
    END
  END mem_in1[27]
  PIN mem_in1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 391.700000 0.600000 391.900000 ;
    END
  END mem_in1[26]
  PIN mem_in1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 391.300000 0.600000 391.500000 ;
    END
  END mem_in1[25]
  PIN mem_in1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 390.900000 0.600000 391.100000 ;
    END
  END mem_in1[24]
  PIN mem_in1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 390.500000 0.600000 390.700000 ;
    END
  END mem_in1[23]
  PIN mem_in1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 390.100000 0.600000 390.300000 ;
    END
  END mem_in1[22]
  PIN mem_in1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.700000 0.600000 389.900000 ;
    END
  END mem_in1[21]
  PIN mem_in1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.300000 0.600000 389.500000 ;
    END
  END mem_in1[20]
  PIN mem_in1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 388.900000 0.600000 389.100000 ;
    END
  END mem_in1[19]
  PIN mem_in1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 388.500000 0.600000 388.700000 ;
    END
  END mem_in1[18]
  PIN mem_in1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 388.100000 0.600000 388.300000 ;
    END
  END mem_in1[17]
  PIN mem_in1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 387.700000 0.600000 387.900000 ;
    END
  END mem_in1[16]
  PIN mem_in1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 387.300000 0.600000 387.500000 ;
    END
  END mem_in1[15]
  PIN mem_in1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.900000 0.600000 387.100000 ;
    END
  END mem_in1[14]
  PIN mem_in1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.500000 0.600000 386.700000 ;
    END
  END mem_in1[13]
  PIN mem_in1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.100000 0.600000 386.300000 ;
    END
  END mem_in1[12]
  PIN mem_in1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 385.700000 0.600000 385.900000 ;
    END
  END mem_in1[11]
  PIN mem_in1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 385.300000 0.600000 385.500000 ;
    END
  END mem_in1[10]
  PIN mem_in1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.900000 0.600000 385.100000 ;
    END
  END mem_in1[9]
  PIN mem_in1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.500000 0.600000 384.700000 ;
    END
  END mem_in1[8]
  PIN mem_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.100000 0.600000 384.300000 ;
    END
  END mem_in1[7]
  PIN mem_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 383.700000 0.600000 383.900000 ;
    END
  END mem_in1[6]
  PIN mem_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 383.300000 0.600000 383.500000 ;
    END
  END mem_in1[5]
  PIN mem_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 382.900000 0.600000 383.100000 ;
    END
  END mem_in1[4]
  PIN mem_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 382.500000 0.600000 382.700000 ;
    END
  END mem_in1[3]
  PIN mem_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 382.100000 0.600000 382.300000 ;
    END
  END mem_in1[2]
  PIN mem_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 381.700000 0.600000 381.900000 ;
    END
  END mem_in1[1]
  PIN mem_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 381.300000 0.600000 381.500000 ;
    END
  END mem_in1[0]
  PIN inst1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[38]
  PIN inst1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[37]
  PIN inst1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[36]
  PIN inst1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[35]
  PIN inst1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[34]
  PIN inst1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[33]
  PIN inst1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[32]
  PIN inst1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[31]
  PIN inst1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[30]
  PIN inst1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst1[29]
  PIN inst1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.300000 0.600000 369.500000 ;
    END
  END inst1[28]
  PIN inst1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 368.900000 0.600000 369.100000 ;
    END
  END inst1[27]
  PIN inst1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 368.500000 0.600000 368.700000 ;
    END
  END inst1[26]
  PIN inst1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 368.100000 0.600000 368.300000 ;
    END
  END inst1[25]
  PIN inst1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 367.700000 0.600000 367.900000 ;
    END
  END inst1[24]
  PIN inst1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 367.300000 0.600000 367.500000 ;
    END
  END inst1[23]
  PIN inst1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 366.900000 0.600000 367.100000 ;
    END
  END inst1[22]
  PIN inst1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 366.500000 0.600000 366.700000 ;
    END
  END inst1[21]
  PIN inst1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 366.100000 0.600000 366.300000 ;
    END
  END inst1[20]
  PIN inst1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 365.700000 0.600000 365.900000 ;
    END
  END inst1[19]
  PIN inst1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 365.300000 0.600000 365.500000 ;
    END
  END inst1[18]
  PIN inst1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.900000 0.600000 365.100000 ;
    END
  END inst1[17]
  PIN inst1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.500000 0.600000 364.700000 ;
    END
  END inst1[16]
  PIN inst1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.100000 0.600000 364.300000 ;
    END
  END inst1[15]
  PIN inst1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 363.700000 0.600000 363.900000 ;
    END
  END inst1[14]
  PIN inst1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 363.300000 0.600000 363.500000 ;
    END
  END inst1[13]
  PIN inst1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 362.900000 0.600000 363.100000 ;
    END
  END inst1[12]
  PIN inst1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 362.500000 0.600000 362.700000 ;
    END
  END inst1[11]
  PIN inst1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 362.100000 0.600000 362.300000 ;
    END
  END inst1[10]
  PIN inst1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 361.700000 0.600000 361.900000 ;
    END
  END inst1[9]
  PIN inst1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 361.300000 0.600000 361.500000 ;
    END
  END inst1[8]
  PIN inst1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 360.900000 0.600000 361.100000 ;
    END
  END inst1[7]
  PIN inst1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 360.500000 0.600000 360.700000 ;
    END
  END inst1[6]
  PIN inst1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 360.100000 0.600000 360.300000 ;
    END
  END inst1[5]
  PIN inst1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 359.700000 0.600000 359.900000 ;
    END
  END inst1[4]
  PIN inst1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 359.300000 0.600000 359.500000 ;
    END
  END inst1[3]
  PIN inst1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 358.900000 0.600000 359.100000 ;
    END
  END inst1[2]
  PIN inst1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 358.500000 0.600000 358.700000 ;
    END
  END inst1[1]
  PIN inst1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 358.100000 0.600000 358.300000 ;
    END
  END inst1[0]
  PIN reset1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 406.900000 0.600000 407.100000 ;
    END
  END reset1
  PIN pmem_out1[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.800000 0.000000 383.000000 0.600000 ;
    END
  END pmem_out1[191]
  PIN pmem_out1[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.400000 0.000000 382.600000 0.600000 ;
    END
  END pmem_out1[190]
  PIN pmem_out1[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.000000 0.000000 382.200000 0.600000 ;
    END
  END pmem_out1[189]
  PIN pmem_out1[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.600000 0.000000 381.800000 0.600000 ;
    END
  END pmem_out1[188]
  PIN pmem_out1[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.200000 0.000000 381.400000 0.600000 ;
    END
  END pmem_out1[187]
  PIN pmem_out1[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.800000 0.000000 381.000000 0.600000 ;
    END
  END pmem_out1[186]
  PIN pmem_out1[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.400000 0.000000 380.600000 0.600000 ;
    END
  END pmem_out1[185]
  PIN pmem_out1[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.000000 0.000000 380.200000 0.600000 ;
    END
  END pmem_out1[184]
  PIN pmem_out1[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.600000 0.000000 379.800000 0.600000 ;
    END
  END pmem_out1[183]
  PIN pmem_out1[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.200000 0.000000 379.400000 0.600000 ;
    END
  END pmem_out1[182]
  PIN pmem_out1[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.800000 0.000000 379.000000 0.600000 ;
    END
  END pmem_out1[181]
  PIN pmem_out1[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.400000 0.000000 378.600000 0.600000 ;
    END
  END pmem_out1[180]
  PIN pmem_out1[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.000000 0.000000 378.200000 0.600000 ;
    END
  END pmem_out1[179]
  PIN pmem_out1[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.600000 0.000000 377.800000 0.600000 ;
    END
  END pmem_out1[178]
  PIN pmem_out1[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.200000 0.000000 377.400000 0.600000 ;
    END
  END pmem_out1[177]
  PIN pmem_out1[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.800000 0.000000 377.000000 0.600000 ;
    END
  END pmem_out1[176]
  PIN pmem_out1[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.400000 0.000000 376.600000 0.600000 ;
    END
  END pmem_out1[175]
  PIN pmem_out1[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.000000 0.000000 376.200000 0.600000 ;
    END
  END pmem_out1[174]
  PIN pmem_out1[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.600000 0.000000 375.800000 0.600000 ;
    END
  END pmem_out1[173]
  PIN pmem_out1[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.200000 0.000000 375.400000 0.600000 ;
    END
  END pmem_out1[172]
  PIN pmem_out1[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.800000 0.000000 375.000000 0.600000 ;
    END
  END pmem_out1[171]
  PIN pmem_out1[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.400000 0.000000 374.600000 0.600000 ;
    END
  END pmem_out1[170]
  PIN pmem_out1[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.000000 0.000000 374.200000 0.600000 ;
    END
  END pmem_out1[169]
  PIN pmem_out1[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.600000 0.000000 373.800000 0.600000 ;
    END
  END pmem_out1[168]
  PIN pmem_out1[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.200000 0.000000 373.400000 0.600000 ;
    END
  END pmem_out1[167]
  PIN pmem_out1[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.800000 0.000000 373.000000 0.600000 ;
    END
  END pmem_out1[166]
  PIN pmem_out1[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.400000 0.000000 372.600000 0.600000 ;
    END
  END pmem_out1[165]
  PIN pmem_out1[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.000000 0.000000 372.200000 0.600000 ;
    END
  END pmem_out1[164]
  PIN pmem_out1[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.600000 0.000000 371.800000 0.600000 ;
    END
  END pmem_out1[163]
  PIN pmem_out1[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.200000 0.000000 371.400000 0.600000 ;
    END
  END pmem_out1[162]
  PIN pmem_out1[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.800000 0.000000 371.000000 0.600000 ;
    END
  END pmem_out1[161]
  PIN pmem_out1[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.400000 0.000000 370.600000 0.600000 ;
    END
  END pmem_out1[160]
  PIN pmem_out1[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.000000 0.000000 370.200000 0.600000 ;
    END
  END pmem_out1[159]
  PIN pmem_out1[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.600000 0.000000 369.800000 0.600000 ;
    END
  END pmem_out1[158]
  PIN pmem_out1[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.200000 0.000000 369.400000 0.600000 ;
    END
  END pmem_out1[157]
  PIN pmem_out1[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.800000 0.000000 369.000000 0.600000 ;
    END
  END pmem_out1[156]
  PIN pmem_out1[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.400000 0.000000 368.600000 0.600000 ;
    END
  END pmem_out1[155]
  PIN pmem_out1[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.000000 0.000000 368.200000 0.600000 ;
    END
  END pmem_out1[154]
  PIN pmem_out1[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.600000 0.000000 367.800000 0.600000 ;
    END
  END pmem_out1[153]
  PIN pmem_out1[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.200000 0.000000 367.400000 0.600000 ;
    END
  END pmem_out1[152]
  PIN pmem_out1[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.800000 0.000000 367.000000 0.600000 ;
    END
  END pmem_out1[151]
  PIN pmem_out1[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.400000 0.000000 366.600000 0.600000 ;
    END
  END pmem_out1[150]
  PIN pmem_out1[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.000000 0.000000 366.200000 0.600000 ;
    END
  END pmem_out1[149]
  PIN pmem_out1[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.600000 0.000000 365.800000 0.600000 ;
    END
  END pmem_out1[148]
  PIN pmem_out1[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.200000 0.000000 365.400000 0.600000 ;
    END
  END pmem_out1[147]
  PIN pmem_out1[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.800000 0.000000 365.000000 0.600000 ;
    END
  END pmem_out1[146]
  PIN pmem_out1[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.400000 0.000000 364.600000 0.600000 ;
    END
  END pmem_out1[145]
  PIN pmem_out1[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.000000 0.000000 364.200000 0.600000 ;
    END
  END pmem_out1[144]
  PIN pmem_out1[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.600000 0.000000 363.800000 0.600000 ;
    END
  END pmem_out1[143]
  PIN pmem_out1[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.200000 0.000000 363.400000 0.600000 ;
    END
  END pmem_out1[142]
  PIN pmem_out1[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.800000 0.000000 363.000000 0.600000 ;
    END
  END pmem_out1[141]
  PIN pmem_out1[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.400000 0.000000 362.600000 0.600000 ;
    END
  END pmem_out1[140]
  PIN pmem_out1[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.000000 0.000000 362.200000 0.600000 ;
    END
  END pmem_out1[139]
  PIN pmem_out1[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.600000 0.000000 361.800000 0.600000 ;
    END
  END pmem_out1[138]
  PIN pmem_out1[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.200000 0.000000 361.400000 0.600000 ;
    END
  END pmem_out1[137]
  PIN pmem_out1[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.800000 0.000000 361.000000 0.600000 ;
    END
  END pmem_out1[136]
  PIN pmem_out1[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.400000 0.000000 360.600000 0.600000 ;
    END
  END pmem_out1[135]
  PIN pmem_out1[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.000000 0.000000 360.200000 0.600000 ;
    END
  END pmem_out1[134]
  PIN pmem_out1[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.600000 0.000000 359.800000 0.600000 ;
    END
  END pmem_out1[133]
  PIN pmem_out1[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.200000 0.000000 359.400000 0.600000 ;
    END
  END pmem_out1[132]
  PIN pmem_out1[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.800000 0.000000 359.000000 0.600000 ;
    END
  END pmem_out1[131]
  PIN pmem_out1[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.400000 0.000000 358.600000 0.600000 ;
    END
  END pmem_out1[130]
  PIN pmem_out1[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.000000 0.000000 358.200000 0.600000 ;
    END
  END pmem_out1[129]
  PIN pmem_out1[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.600000 0.000000 357.800000 0.600000 ;
    END
  END pmem_out1[128]
  PIN pmem_out1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.200000 0.000000 357.400000 0.600000 ;
    END
  END pmem_out1[127]
  PIN pmem_out1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.800000 0.000000 357.000000 0.600000 ;
    END
  END pmem_out1[126]
  PIN pmem_out1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.400000 0.000000 356.600000 0.600000 ;
    END
  END pmem_out1[125]
  PIN pmem_out1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.000000 0.000000 356.200000 0.600000 ;
    END
  END pmem_out1[124]
  PIN pmem_out1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.600000 0.000000 355.800000 0.600000 ;
    END
  END pmem_out1[123]
  PIN pmem_out1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.200000 0.000000 355.400000 0.600000 ;
    END
  END pmem_out1[122]
  PIN pmem_out1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.800000 0.000000 355.000000 0.600000 ;
    END
  END pmem_out1[121]
  PIN pmem_out1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.400000 0.000000 354.600000 0.600000 ;
    END
  END pmem_out1[120]
  PIN pmem_out1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.000000 0.000000 354.200000 0.600000 ;
    END
  END pmem_out1[119]
  PIN pmem_out1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.600000 0.000000 353.800000 0.600000 ;
    END
  END pmem_out1[118]
  PIN pmem_out1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.200000 0.000000 353.400000 0.600000 ;
    END
  END pmem_out1[117]
  PIN pmem_out1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.800000 0.000000 353.000000 0.600000 ;
    END
  END pmem_out1[116]
  PIN pmem_out1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.400000 0.000000 352.600000 0.600000 ;
    END
  END pmem_out1[115]
  PIN pmem_out1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.000000 0.000000 352.200000 0.600000 ;
    END
  END pmem_out1[114]
  PIN pmem_out1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.600000 0.000000 351.800000 0.600000 ;
    END
  END pmem_out1[113]
  PIN pmem_out1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.200000 0.000000 351.400000 0.600000 ;
    END
  END pmem_out1[112]
  PIN pmem_out1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.800000 0.000000 351.000000 0.600000 ;
    END
  END pmem_out1[111]
  PIN pmem_out1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.400000 0.000000 350.600000 0.600000 ;
    END
  END pmem_out1[110]
  PIN pmem_out1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.000000 0.000000 350.200000 0.600000 ;
    END
  END pmem_out1[109]
  PIN pmem_out1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.600000 0.000000 349.800000 0.600000 ;
    END
  END pmem_out1[108]
  PIN pmem_out1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.200000 0.000000 349.400000 0.600000 ;
    END
  END pmem_out1[107]
  PIN pmem_out1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.800000 0.000000 349.000000 0.600000 ;
    END
  END pmem_out1[106]
  PIN pmem_out1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.400000 0.000000 348.600000 0.600000 ;
    END
  END pmem_out1[105]
  PIN pmem_out1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.000000 0.000000 348.200000 0.600000 ;
    END
  END pmem_out1[104]
  PIN pmem_out1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.600000 0.000000 347.800000 0.600000 ;
    END
  END pmem_out1[103]
  PIN pmem_out1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.200000 0.000000 347.400000 0.600000 ;
    END
  END pmem_out1[102]
  PIN pmem_out1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.800000 0.000000 347.000000 0.600000 ;
    END
  END pmem_out1[101]
  PIN pmem_out1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.400000 0.000000 346.600000 0.600000 ;
    END
  END pmem_out1[100]
  PIN pmem_out1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.000000 0.000000 346.200000 0.600000 ;
    END
  END pmem_out1[99]
  PIN pmem_out1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.600000 0.000000 345.800000 0.600000 ;
    END
  END pmem_out1[98]
  PIN pmem_out1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.200000 0.000000 345.400000 0.600000 ;
    END
  END pmem_out1[97]
  PIN pmem_out1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.800000 0.000000 345.000000 0.600000 ;
    END
  END pmem_out1[96]
  PIN pmem_out1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.400000 0.000000 344.600000 0.600000 ;
    END
  END pmem_out1[95]
  PIN pmem_out1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.000000 0.000000 344.200000 0.600000 ;
    END
  END pmem_out1[94]
  PIN pmem_out1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.600000 0.000000 343.800000 0.600000 ;
    END
  END pmem_out1[93]
  PIN pmem_out1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.200000 0.000000 343.400000 0.600000 ;
    END
  END pmem_out1[92]
  PIN pmem_out1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.800000 0.000000 343.000000 0.600000 ;
    END
  END pmem_out1[91]
  PIN pmem_out1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.400000 0.000000 342.600000 0.600000 ;
    END
  END pmem_out1[90]
  PIN pmem_out1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.000000 0.000000 342.200000 0.600000 ;
    END
  END pmem_out1[89]
  PIN pmem_out1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.600000 0.000000 341.800000 0.600000 ;
    END
  END pmem_out1[88]
  PIN pmem_out1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.200000 0.000000 341.400000 0.600000 ;
    END
  END pmem_out1[87]
  PIN pmem_out1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.800000 0.000000 341.000000 0.600000 ;
    END
  END pmem_out1[86]
  PIN pmem_out1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.400000 0.000000 340.600000 0.600000 ;
    END
  END pmem_out1[85]
  PIN pmem_out1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.000000 0.000000 340.200000 0.600000 ;
    END
  END pmem_out1[84]
  PIN pmem_out1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.600000 0.000000 339.800000 0.600000 ;
    END
  END pmem_out1[83]
  PIN pmem_out1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.200000 0.000000 339.400000 0.600000 ;
    END
  END pmem_out1[82]
  PIN pmem_out1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.800000 0.000000 339.000000 0.600000 ;
    END
  END pmem_out1[81]
  PIN pmem_out1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.400000 0.000000 338.600000 0.600000 ;
    END
  END pmem_out1[80]
  PIN pmem_out1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.000000 0.000000 338.200000 0.600000 ;
    END
  END pmem_out1[79]
  PIN pmem_out1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.600000 0.000000 337.800000 0.600000 ;
    END
  END pmem_out1[78]
  PIN pmem_out1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.200000 0.000000 337.400000 0.600000 ;
    END
  END pmem_out1[77]
  PIN pmem_out1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.800000 0.000000 337.000000 0.600000 ;
    END
  END pmem_out1[76]
  PIN pmem_out1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.400000 0.000000 336.600000 0.600000 ;
    END
  END pmem_out1[75]
  PIN pmem_out1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.000000 0.000000 336.200000 0.600000 ;
    END
  END pmem_out1[74]
  PIN pmem_out1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.600000 0.000000 335.800000 0.600000 ;
    END
  END pmem_out1[73]
  PIN pmem_out1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.200000 0.000000 335.400000 0.600000 ;
    END
  END pmem_out1[72]
  PIN pmem_out1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.800000 0.000000 335.000000 0.600000 ;
    END
  END pmem_out1[71]
  PIN pmem_out1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.400000 0.000000 334.600000 0.600000 ;
    END
  END pmem_out1[70]
  PIN pmem_out1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.000000 0.000000 334.200000 0.600000 ;
    END
  END pmem_out1[69]
  PIN pmem_out1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.600000 0.000000 333.800000 0.600000 ;
    END
  END pmem_out1[68]
  PIN pmem_out1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.200000 0.000000 333.400000 0.600000 ;
    END
  END pmem_out1[67]
  PIN pmem_out1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.800000 0.000000 333.000000 0.600000 ;
    END
  END pmem_out1[66]
  PIN pmem_out1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.400000 0.000000 332.600000 0.600000 ;
    END
  END pmem_out1[65]
  PIN pmem_out1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.000000 0.000000 332.200000 0.600000 ;
    END
  END pmem_out1[64]
  PIN pmem_out1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.600000 0.000000 331.800000 0.600000 ;
    END
  END pmem_out1[63]
  PIN pmem_out1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.200000 0.000000 331.400000 0.600000 ;
    END
  END pmem_out1[62]
  PIN pmem_out1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.800000 0.000000 331.000000 0.600000 ;
    END
  END pmem_out1[61]
  PIN pmem_out1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.400000 0.000000 330.600000 0.600000 ;
    END
  END pmem_out1[60]
  PIN pmem_out1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.000000 0.000000 330.200000 0.600000 ;
    END
  END pmem_out1[59]
  PIN pmem_out1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.600000 0.000000 329.800000 0.600000 ;
    END
  END pmem_out1[58]
  PIN pmem_out1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.200000 0.000000 329.400000 0.600000 ;
    END
  END pmem_out1[57]
  PIN pmem_out1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.800000 0.000000 329.000000 0.600000 ;
    END
  END pmem_out1[56]
  PIN pmem_out1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.400000 0.000000 328.600000 0.600000 ;
    END
  END pmem_out1[55]
  PIN pmem_out1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.000000 0.000000 328.200000 0.600000 ;
    END
  END pmem_out1[54]
  PIN pmem_out1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.600000 0.000000 327.800000 0.600000 ;
    END
  END pmem_out1[53]
  PIN pmem_out1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.200000 0.000000 327.400000 0.600000 ;
    END
  END pmem_out1[52]
  PIN pmem_out1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.800000 0.000000 327.000000 0.600000 ;
    END
  END pmem_out1[51]
  PIN pmem_out1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.400000 0.000000 326.600000 0.600000 ;
    END
  END pmem_out1[50]
  PIN pmem_out1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.000000 0.000000 326.200000 0.600000 ;
    END
  END pmem_out1[49]
  PIN pmem_out1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.600000 0.000000 325.800000 0.600000 ;
    END
  END pmem_out1[48]
  PIN pmem_out1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.200000 0.000000 325.400000 0.600000 ;
    END
  END pmem_out1[47]
  PIN pmem_out1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.800000 0.000000 325.000000 0.600000 ;
    END
  END pmem_out1[46]
  PIN pmem_out1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.400000 0.000000 324.600000 0.600000 ;
    END
  END pmem_out1[45]
  PIN pmem_out1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.000000 0.000000 324.200000 0.600000 ;
    END
  END pmem_out1[44]
  PIN pmem_out1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.600000 0.000000 323.800000 0.600000 ;
    END
  END pmem_out1[43]
  PIN pmem_out1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.200000 0.000000 323.400000 0.600000 ;
    END
  END pmem_out1[42]
  PIN pmem_out1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.800000 0.000000 323.000000 0.600000 ;
    END
  END pmem_out1[41]
  PIN pmem_out1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.400000 0.000000 322.600000 0.600000 ;
    END
  END pmem_out1[40]
  PIN pmem_out1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.000000 0.000000 322.200000 0.600000 ;
    END
  END pmem_out1[39]
  PIN pmem_out1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.600000 0.000000 321.800000 0.600000 ;
    END
  END pmem_out1[38]
  PIN pmem_out1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.200000 0.000000 321.400000 0.600000 ;
    END
  END pmem_out1[37]
  PIN pmem_out1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.800000 0.000000 321.000000 0.600000 ;
    END
  END pmem_out1[36]
  PIN pmem_out1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.400000 0.000000 320.600000 0.600000 ;
    END
  END pmem_out1[35]
  PIN pmem_out1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.000000 0.000000 320.200000 0.600000 ;
    END
  END pmem_out1[34]
  PIN pmem_out1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.600000 0.000000 319.800000 0.600000 ;
    END
  END pmem_out1[33]
  PIN pmem_out1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.200000 0.000000 319.400000 0.600000 ;
    END
  END pmem_out1[32]
  PIN pmem_out1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.800000 0.000000 319.000000 0.600000 ;
    END
  END pmem_out1[31]
  PIN pmem_out1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.400000 0.000000 318.600000 0.600000 ;
    END
  END pmem_out1[30]
  PIN pmem_out1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.000000 0.000000 318.200000 0.600000 ;
    END
  END pmem_out1[29]
  PIN pmem_out1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.600000 0.000000 317.800000 0.600000 ;
    END
  END pmem_out1[28]
  PIN pmem_out1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.200000 0.000000 317.400000 0.600000 ;
    END
  END pmem_out1[27]
  PIN pmem_out1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.800000 0.000000 317.000000 0.600000 ;
    END
  END pmem_out1[26]
  PIN pmem_out1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.400000 0.000000 316.600000 0.600000 ;
    END
  END pmem_out1[25]
  PIN pmem_out1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.000000 0.000000 316.200000 0.600000 ;
    END
  END pmem_out1[24]
  PIN pmem_out1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.600000 0.000000 315.800000 0.600000 ;
    END
  END pmem_out1[23]
  PIN pmem_out1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.200000 0.000000 315.400000 0.600000 ;
    END
  END pmem_out1[22]
  PIN pmem_out1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.800000 0.000000 315.000000 0.600000 ;
    END
  END pmem_out1[21]
  PIN pmem_out1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.400000 0.000000 314.600000 0.600000 ;
    END
  END pmem_out1[20]
  PIN pmem_out1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.000000 0.000000 314.200000 0.600000 ;
    END
  END pmem_out1[19]
  PIN pmem_out1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.600000 0.000000 313.800000 0.600000 ;
    END
  END pmem_out1[18]
  PIN pmem_out1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.200000 0.000000 313.400000 0.600000 ;
    END
  END pmem_out1[17]
  PIN pmem_out1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.800000 0.000000 313.000000 0.600000 ;
    END
  END pmem_out1[16]
  PIN pmem_out1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.400000 0.000000 312.600000 0.600000 ;
    END
  END pmem_out1[15]
  PIN pmem_out1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.000000 0.000000 312.200000 0.600000 ;
    END
  END pmem_out1[14]
  PIN pmem_out1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.600000 0.000000 311.800000 0.600000 ;
    END
  END pmem_out1[13]
  PIN pmem_out1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.200000 0.000000 311.400000 0.600000 ;
    END
  END pmem_out1[12]
  PIN pmem_out1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.800000 0.000000 311.000000 0.600000 ;
    END
  END pmem_out1[11]
  PIN pmem_out1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.400000 0.000000 310.600000 0.600000 ;
    END
  END pmem_out1[10]
  PIN pmem_out1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.000000 0.000000 310.200000 0.600000 ;
    END
  END pmem_out1[9]
  PIN pmem_out1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.600000 0.000000 309.800000 0.600000 ;
    END
  END pmem_out1[8]
  PIN pmem_out1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.200000 0.000000 309.400000 0.600000 ;
    END
  END pmem_out1[7]
  PIN pmem_out1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.800000 0.000000 309.000000 0.600000 ;
    END
  END pmem_out1[6]
  PIN pmem_out1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.400000 0.000000 308.600000 0.600000 ;
    END
  END pmem_out1[5]
  PIN pmem_out1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.000000 0.000000 308.200000 0.600000 ;
    END
  END pmem_out1[4]
  PIN pmem_out1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.600000 0.000000 307.800000 0.600000 ;
    END
  END pmem_out1[3]
  PIN pmem_out1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.200000 0.000000 307.400000 0.600000 ;
    END
  END pmem_out1[2]
  PIN pmem_out1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.800000 0.000000 307.000000 0.600000 ;
    END
  END pmem_out1[1]
  PIN pmem_out1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.400000 0.000000 306.600000 0.600000 ;
    END
  END pmem_out1[0]
  PIN mem_in2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 406.500000 0.600000 406.700000 ;
    END
  END mem_in2[31]
  PIN mem_in2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 406.100000 0.600000 406.300000 ;
    END
  END mem_in2[30]
  PIN mem_in2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 405.700000 0.600000 405.900000 ;
    END
  END mem_in2[29]
  PIN mem_in2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 405.300000 0.600000 405.500000 ;
    END
  END mem_in2[28]
  PIN mem_in2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.900000 0.600000 405.100000 ;
    END
  END mem_in2[27]
  PIN mem_in2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.500000 0.600000 404.700000 ;
    END
  END mem_in2[26]
  PIN mem_in2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.100000 0.600000 404.300000 ;
    END
  END mem_in2[25]
  PIN mem_in2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 403.700000 0.600000 403.900000 ;
    END
  END mem_in2[24]
  PIN mem_in2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 403.300000 0.600000 403.500000 ;
    END
  END mem_in2[23]
  PIN mem_in2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 402.900000 0.600000 403.100000 ;
    END
  END mem_in2[22]
  PIN mem_in2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 402.500000 0.600000 402.700000 ;
    END
  END mem_in2[21]
  PIN mem_in2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 402.100000 0.600000 402.300000 ;
    END
  END mem_in2[20]
  PIN mem_in2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 401.700000 0.600000 401.900000 ;
    END
  END mem_in2[19]
  PIN mem_in2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 401.300000 0.600000 401.500000 ;
    END
  END mem_in2[18]
  PIN mem_in2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 400.900000 0.600000 401.100000 ;
    END
  END mem_in2[17]
  PIN mem_in2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 400.500000 0.600000 400.700000 ;
    END
  END mem_in2[16]
  PIN mem_in2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 400.100000 0.600000 400.300000 ;
    END
  END mem_in2[15]
  PIN mem_in2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 399.700000 0.600000 399.900000 ;
    END
  END mem_in2[14]
  PIN mem_in2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 399.300000 0.600000 399.500000 ;
    END
  END mem_in2[13]
  PIN mem_in2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.900000 0.600000 399.100000 ;
    END
  END mem_in2[12]
  PIN mem_in2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.500000 0.600000 398.700000 ;
    END
  END mem_in2[11]
  PIN mem_in2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.100000 0.600000 398.300000 ;
    END
  END mem_in2[10]
  PIN mem_in2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 397.700000 0.600000 397.900000 ;
    END
  END mem_in2[9]
  PIN mem_in2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 397.300000 0.600000 397.500000 ;
    END
  END mem_in2[8]
  PIN mem_in2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 396.900000 0.600000 397.100000 ;
    END
  END mem_in2[7]
  PIN mem_in2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 396.500000 0.600000 396.700000 ;
    END
  END mem_in2[6]
  PIN mem_in2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 396.100000 0.600000 396.300000 ;
    END
  END mem_in2[5]
  PIN mem_in2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 395.700000 0.600000 395.900000 ;
    END
  END mem_in2[4]
  PIN mem_in2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 395.300000 0.600000 395.500000 ;
    END
  END mem_in2[3]
  PIN mem_in2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.900000 0.600000 395.100000 ;
    END
  END mem_in2[2]
  PIN mem_in2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.500000 0.600000 394.700000 ;
    END
  END mem_in2[1]
  PIN mem_in2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.100000 0.600000 394.300000 ;
    END
  END mem_in2[0]
  PIN inst2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[38]
  PIN inst2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[37]
  PIN inst2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[36]
  PIN inst2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[35]
  PIN inst2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[34]
  PIN inst2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[33]
  PIN inst2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[32]
  PIN inst2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[31]
  PIN inst2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[30]
  PIN inst2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END inst2[29]
  PIN inst2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 380.900000 0.600000 381.100000 ;
    END
  END inst2[28]
  PIN inst2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 380.500000 0.600000 380.700000 ;
    END
  END inst2[27]
  PIN inst2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 380.100000 0.600000 380.300000 ;
    END
  END inst2[26]
  PIN inst2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 379.700000 0.600000 379.900000 ;
    END
  END inst2[25]
  PIN inst2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 379.300000 0.600000 379.500000 ;
    END
  END inst2[24]
  PIN inst2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 378.900000 0.600000 379.100000 ;
    END
  END inst2[23]
  PIN inst2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 378.500000 0.600000 378.700000 ;
    END
  END inst2[22]
  PIN inst2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 378.100000 0.600000 378.300000 ;
    END
  END inst2[21]
  PIN inst2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 377.700000 0.600000 377.900000 ;
    END
  END inst2[20]
  PIN inst2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 377.300000 0.600000 377.500000 ;
    END
  END inst2[19]
  PIN inst2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 376.900000 0.600000 377.100000 ;
    END
  END inst2[18]
  PIN inst2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 376.500000 0.600000 376.700000 ;
    END
  END inst2[17]
  PIN inst2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 376.100000 0.600000 376.300000 ;
    END
  END inst2[16]
  PIN inst2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 375.700000 0.600000 375.900000 ;
    END
  END inst2[15]
  PIN inst2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 375.300000 0.600000 375.500000 ;
    END
  END inst2[14]
  PIN inst2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 374.900000 0.600000 375.100000 ;
    END
  END inst2[13]
  PIN inst2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 374.500000 0.600000 374.700000 ;
    END
  END inst2[12]
  PIN inst2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 374.100000 0.600000 374.300000 ;
    END
  END inst2[11]
  PIN inst2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 373.700000 0.600000 373.900000 ;
    END
  END inst2[10]
  PIN inst2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 373.300000 0.600000 373.500000 ;
    END
  END inst2[9]
  PIN inst2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 372.900000 0.600000 373.100000 ;
    END
  END inst2[8]
  PIN inst2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 372.500000 0.600000 372.700000 ;
    END
  END inst2[7]
  PIN inst2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 372.100000 0.600000 372.300000 ;
    END
  END inst2[6]
  PIN inst2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 371.700000 0.600000 371.900000 ;
    END
  END inst2[5]
  PIN inst2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 371.300000 0.600000 371.500000 ;
    END
  END inst2[4]
  PIN inst2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 370.900000 0.600000 371.100000 ;
    END
  END inst2[3]
  PIN inst2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 370.500000 0.600000 370.700000 ;
    END
  END inst2[2]
  PIN inst2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 370.100000 0.600000 370.300000 ;
    END
  END inst2[1]
  PIN inst2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.700000 0.600000 369.900000 ;
    END
  END inst2[0]
  PIN reset2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 407.300000 0.600000 407.500000 ;
    END
  END reset2
  PIN pmem_out2[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.600000 0.000000 459.800000 0.600000 ;
    END
  END pmem_out2[191]
  PIN pmem_out2[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.200000 0.000000 459.400000 0.600000 ;
    END
  END pmem_out2[190]
  PIN pmem_out2[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.800000 0.000000 459.000000 0.600000 ;
    END
  END pmem_out2[189]
  PIN pmem_out2[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.400000 0.000000 458.600000 0.600000 ;
    END
  END pmem_out2[188]
  PIN pmem_out2[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.000000 0.000000 458.200000 0.600000 ;
    END
  END pmem_out2[187]
  PIN pmem_out2[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.600000 0.000000 457.800000 0.600000 ;
    END
  END pmem_out2[186]
  PIN pmem_out2[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.200000 0.000000 457.400000 0.600000 ;
    END
  END pmem_out2[185]
  PIN pmem_out2[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.800000 0.000000 457.000000 0.600000 ;
    END
  END pmem_out2[184]
  PIN pmem_out2[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.400000 0.000000 456.600000 0.600000 ;
    END
  END pmem_out2[183]
  PIN pmem_out2[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.000000 0.000000 456.200000 0.600000 ;
    END
  END pmem_out2[182]
  PIN pmem_out2[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.600000 0.000000 455.800000 0.600000 ;
    END
  END pmem_out2[181]
  PIN pmem_out2[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.200000 0.000000 455.400000 0.600000 ;
    END
  END pmem_out2[180]
  PIN pmem_out2[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.800000 0.000000 455.000000 0.600000 ;
    END
  END pmem_out2[179]
  PIN pmem_out2[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.400000 0.000000 454.600000 0.600000 ;
    END
  END pmem_out2[178]
  PIN pmem_out2[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.000000 0.000000 454.200000 0.600000 ;
    END
  END pmem_out2[177]
  PIN pmem_out2[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.600000 0.000000 453.800000 0.600000 ;
    END
  END pmem_out2[176]
  PIN pmem_out2[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.200000 0.000000 453.400000 0.600000 ;
    END
  END pmem_out2[175]
  PIN pmem_out2[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.800000 0.000000 453.000000 0.600000 ;
    END
  END pmem_out2[174]
  PIN pmem_out2[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.400000 0.000000 452.600000 0.600000 ;
    END
  END pmem_out2[173]
  PIN pmem_out2[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.000000 0.000000 452.200000 0.600000 ;
    END
  END pmem_out2[172]
  PIN pmem_out2[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.600000 0.000000 451.800000 0.600000 ;
    END
  END pmem_out2[171]
  PIN pmem_out2[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.200000 0.000000 451.400000 0.600000 ;
    END
  END pmem_out2[170]
  PIN pmem_out2[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.800000 0.000000 451.000000 0.600000 ;
    END
  END pmem_out2[169]
  PIN pmem_out2[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.400000 0.000000 450.600000 0.600000 ;
    END
  END pmem_out2[168]
  PIN pmem_out2[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.000000 0.000000 450.200000 0.600000 ;
    END
  END pmem_out2[167]
  PIN pmem_out2[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.600000 0.000000 449.800000 0.600000 ;
    END
  END pmem_out2[166]
  PIN pmem_out2[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.200000 0.000000 449.400000 0.600000 ;
    END
  END pmem_out2[165]
  PIN pmem_out2[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.800000 0.000000 449.000000 0.600000 ;
    END
  END pmem_out2[164]
  PIN pmem_out2[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.400000 0.000000 448.600000 0.600000 ;
    END
  END pmem_out2[163]
  PIN pmem_out2[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.000000 0.000000 448.200000 0.600000 ;
    END
  END pmem_out2[162]
  PIN pmem_out2[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.600000 0.000000 447.800000 0.600000 ;
    END
  END pmem_out2[161]
  PIN pmem_out2[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.200000 0.000000 447.400000 0.600000 ;
    END
  END pmem_out2[160]
  PIN pmem_out2[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.800000 0.000000 447.000000 0.600000 ;
    END
  END pmem_out2[159]
  PIN pmem_out2[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.400000 0.000000 446.600000 0.600000 ;
    END
  END pmem_out2[158]
  PIN pmem_out2[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.000000 0.000000 446.200000 0.600000 ;
    END
  END pmem_out2[157]
  PIN pmem_out2[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.600000 0.000000 445.800000 0.600000 ;
    END
  END pmem_out2[156]
  PIN pmem_out2[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.200000 0.000000 445.400000 0.600000 ;
    END
  END pmem_out2[155]
  PIN pmem_out2[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.800000 0.000000 445.000000 0.600000 ;
    END
  END pmem_out2[154]
  PIN pmem_out2[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.400000 0.000000 444.600000 0.600000 ;
    END
  END pmem_out2[153]
  PIN pmem_out2[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.000000 0.000000 444.200000 0.600000 ;
    END
  END pmem_out2[152]
  PIN pmem_out2[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.600000 0.000000 443.800000 0.600000 ;
    END
  END pmem_out2[151]
  PIN pmem_out2[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.200000 0.000000 443.400000 0.600000 ;
    END
  END pmem_out2[150]
  PIN pmem_out2[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.800000 0.000000 443.000000 0.600000 ;
    END
  END pmem_out2[149]
  PIN pmem_out2[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.400000 0.000000 442.600000 0.600000 ;
    END
  END pmem_out2[148]
  PIN pmem_out2[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.000000 0.000000 442.200000 0.600000 ;
    END
  END pmem_out2[147]
  PIN pmem_out2[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.600000 0.000000 441.800000 0.600000 ;
    END
  END pmem_out2[146]
  PIN pmem_out2[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.200000 0.000000 441.400000 0.600000 ;
    END
  END pmem_out2[145]
  PIN pmem_out2[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.800000 0.000000 441.000000 0.600000 ;
    END
  END pmem_out2[144]
  PIN pmem_out2[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.400000 0.000000 440.600000 0.600000 ;
    END
  END pmem_out2[143]
  PIN pmem_out2[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.000000 0.000000 440.200000 0.600000 ;
    END
  END pmem_out2[142]
  PIN pmem_out2[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.600000 0.000000 439.800000 0.600000 ;
    END
  END pmem_out2[141]
  PIN pmem_out2[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.200000 0.000000 439.400000 0.600000 ;
    END
  END pmem_out2[140]
  PIN pmem_out2[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.800000 0.000000 439.000000 0.600000 ;
    END
  END pmem_out2[139]
  PIN pmem_out2[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.400000 0.000000 438.600000 0.600000 ;
    END
  END pmem_out2[138]
  PIN pmem_out2[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.000000 0.000000 438.200000 0.600000 ;
    END
  END pmem_out2[137]
  PIN pmem_out2[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.600000 0.000000 437.800000 0.600000 ;
    END
  END pmem_out2[136]
  PIN pmem_out2[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.200000 0.000000 437.400000 0.600000 ;
    END
  END pmem_out2[135]
  PIN pmem_out2[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.800000 0.000000 437.000000 0.600000 ;
    END
  END pmem_out2[134]
  PIN pmem_out2[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.400000 0.000000 436.600000 0.600000 ;
    END
  END pmem_out2[133]
  PIN pmem_out2[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.000000 0.000000 436.200000 0.600000 ;
    END
  END pmem_out2[132]
  PIN pmem_out2[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.600000 0.000000 435.800000 0.600000 ;
    END
  END pmem_out2[131]
  PIN pmem_out2[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.200000 0.000000 435.400000 0.600000 ;
    END
  END pmem_out2[130]
  PIN pmem_out2[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.800000 0.000000 435.000000 0.600000 ;
    END
  END pmem_out2[129]
  PIN pmem_out2[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.400000 0.000000 434.600000 0.600000 ;
    END
  END pmem_out2[128]
  PIN pmem_out2[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.000000 0.000000 434.200000 0.600000 ;
    END
  END pmem_out2[127]
  PIN pmem_out2[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.600000 0.000000 433.800000 0.600000 ;
    END
  END pmem_out2[126]
  PIN pmem_out2[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.200000 0.000000 433.400000 0.600000 ;
    END
  END pmem_out2[125]
  PIN pmem_out2[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.800000 0.000000 433.000000 0.600000 ;
    END
  END pmem_out2[124]
  PIN pmem_out2[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.400000 0.000000 432.600000 0.600000 ;
    END
  END pmem_out2[123]
  PIN pmem_out2[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.000000 0.000000 432.200000 0.600000 ;
    END
  END pmem_out2[122]
  PIN pmem_out2[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.600000 0.000000 431.800000 0.600000 ;
    END
  END pmem_out2[121]
  PIN pmem_out2[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.200000 0.000000 431.400000 0.600000 ;
    END
  END pmem_out2[120]
  PIN pmem_out2[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.800000 0.000000 431.000000 0.600000 ;
    END
  END pmem_out2[119]
  PIN pmem_out2[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.400000 0.000000 430.600000 0.600000 ;
    END
  END pmem_out2[118]
  PIN pmem_out2[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.000000 0.000000 430.200000 0.600000 ;
    END
  END pmem_out2[117]
  PIN pmem_out2[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.600000 0.000000 429.800000 0.600000 ;
    END
  END pmem_out2[116]
  PIN pmem_out2[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.200000 0.000000 429.400000 0.600000 ;
    END
  END pmem_out2[115]
  PIN pmem_out2[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.800000 0.000000 429.000000 0.600000 ;
    END
  END pmem_out2[114]
  PIN pmem_out2[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.400000 0.000000 428.600000 0.600000 ;
    END
  END pmem_out2[113]
  PIN pmem_out2[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.000000 0.000000 428.200000 0.600000 ;
    END
  END pmem_out2[112]
  PIN pmem_out2[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.600000 0.000000 427.800000 0.600000 ;
    END
  END pmem_out2[111]
  PIN pmem_out2[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.200000 0.000000 427.400000 0.600000 ;
    END
  END pmem_out2[110]
  PIN pmem_out2[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.800000 0.000000 427.000000 0.600000 ;
    END
  END pmem_out2[109]
  PIN pmem_out2[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.400000 0.000000 426.600000 0.600000 ;
    END
  END pmem_out2[108]
  PIN pmem_out2[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.000000 0.000000 426.200000 0.600000 ;
    END
  END pmem_out2[107]
  PIN pmem_out2[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.600000 0.000000 425.800000 0.600000 ;
    END
  END pmem_out2[106]
  PIN pmem_out2[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.200000 0.000000 425.400000 0.600000 ;
    END
  END pmem_out2[105]
  PIN pmem_out2[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.800000 0.000000 425.000000 0.600000 ;
    END
  END pmem_out2[104]
  PIN pmem_out2[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.400000 0.000000 424.600000 0.600000 ;
    END
  END pmem_out2[103]
  PIN pmem_out2[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.000000 0.000000 424.200000 0.600000 ;
    END
  END pmem_out2[102]
  PIN pmem_out2[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.600000 0.000000 423.800000 0.600000 ;
    END
  END pmem_out2[101]
  PIN pmem_out2[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.200000 0.000000 423.400000 0.600000 ;
    END
  END pmem_out2[100]
  PIN pmem_out2[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.800000 0.000000 423.000000 0.600000 ;
    END
  END pmem_out2[99]
  PIN pmem_out2[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.400000 0.000000 422.600000 0.600000 ;
    END
  END pmem_out2[98]
  PIN pmem_out2[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.000000 0.000000 422.200000 0.600000 ;
    END
  END pmem_out2[97]
  PIN pmem_out2[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.600000 0.000000 421.800000 0.600000 ;
    END
  END pmem_out2[96]
  PIN pmem_out2[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.200000 0.000000 421.400000 0.600000 ;
    END
  END pmem_out2[95]
  PIN pmem_out2[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.800000 0.000000 421.000000 0.600000 ;
    END
  END pmem_out2[94]
  PIN pmem_out2[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.400000 0.000000 420.600000 0.600000 ;
    END
  END pmem_out2[93]
  PIN pmem_out2[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.000000 0.000000 420.200000 0.600000 ;
    END
  END pmem_out2[92]
  PIN pmem_out2[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.600000 0.000000 419.800000 0.600000 ;
    END
  END pmem_out2[91]
  PIN pmem_out2[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.200000 0.000000 419.400000 0.600000 ;
    END
  END pmem_out2[90]
  PIN pmem_out2[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.800000 0.000000 419.000000 0.600000 ;
    END
  END pmem_out2[89]
  PIN pmem_out2[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.400000 0.000000 418.600000 0.600000 ;
    END
  END pmem_out2[88]
  PIN pmem_out2[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.000000 0.000000 418.200000 0.600000 ;
    END
  END pmem_out2[87]
  PIN pmem_out2[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.600000 0.000000 417.800000 0.600000 ;
    END
  END pmem_out2[86]
  PIN pmem_out2[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.200000 0.000000 417.400000 0.600000 ;
    END
  END pmem_out2[85]
  PIN pmem_out2[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.800000 0.000000 417.000000 0.600000 ;
    END
  END pmem_out2[84]
  PIN pmem_out2[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.400000 0.000000 416.600000 0.600000 ;
    END
  END pmem_out2[83]
  PIN pmem_out2[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.000000 0.000000 416.200000 0.600000 ;
    END
  END pmem_out2[82]
  PIN pmem_out2[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.600000 0.000000 415.800000 0.600000 ;
    END
  END pmem_out2[81]
  PIN pmem_out2[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.200000 0.000000 415.400000 0.600000 ;
    END
  END pmem_out2[80]
  PIN pmem_out2[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.800000 0.000000 415.000000 0.600000 ;
    END
  END pmem_out2[79]
  PIN pmem_out2[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.400000 0.000000 414.600000 0.600000 ;
    END
  END pmem_out2[78]
  PIN pmem_out2[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.000000 0.000000 414.200000 0.600000 ;
    END
  END pmem_out2[77]
  PIN pmem_out2[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.600000 0.000000 413.800000 0.600000 ;
    END
  END pmem_out2[76]
  PIN pmem_out2[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.200000 0.000000 413.400000 0.600000 ;
    END
  END pmem_out2[75]
  PIN pmem_out2[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.800000 0.000000 413.000000 0.600000 ;
    END
  END pmem_out2[74]
  PIN pmem_out2[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.400000 0.000000 412.600000 0.600000 ;
    END
  END pmem_out2[73]
  PIN pmem_out2[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.000000 0.000000 412.200000 0.600000 ;
    END
  END pmem_out2[72]
  PIN pmem_out2[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.600000 0.000000 411.800000 0.600000 ;
    END
  END pmem_out2[71]
  PIN pmem_out2[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.200000 0.000000 411.400000 0.600000 ;
    END
  END pmem_out2[70]
  PIN pmem_out2[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.800000 0.000000 411.000000 0.600000 ;
    END
  END pmem_out2[69]
  PIN pmem_out2[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.400000 0.000000 410.600000 0.600000 ;
    END
  END pmem_out2[68]
  PIN pmem_out2[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.000000 0.000000 410.200000 0.600000 ;
    END
  END pmem_out2[67]
  PIN pmem_out2[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.600000 0.000000 409.800000 0.600000 ;
    END
  END pmem_out2[66]
  PIN pmem_out2[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.200000 0.000000 409.400000 0.600000 ;
    END
  END pmem_out2[65]
  PIN pmem_out2[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.800000 0.000000 409.000000 0.600000 ;
    END
  END pmem_out2[64]
  PIN pmem_out2[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.400000 0.000000 408.600000 0.600000 ;
    END
  END pmem_out2[63]
  PIN pmem_out2[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.000000 0.000000 408.200000 0.600000 ;
    END
  END pmem_out2[62]
  PIN pmem_out2[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.600000 0.000000 407.800000 0.600000 ;
    END
  END pmem_out2[61]
  PIN pmem_out2[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.200000 0.000000 407.400000 0.600000 ;
    END
  END pmem_out2[60]
  PIN pmem_out2[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.800000 0.000000 407.000000 0.600000 ;
    END
  END pmem_out2[59]
  PIN pmem_out2[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.400000 0.000000 406.600000 0.600000 ;
    END
  END pmem_out2[58]
  PIN pmem_out2[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.000000 0.000000 406.200000 0.600000 ;
    END
  END pmem_out2[57]
  PIN pmem_out2[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.600000 0.000000 405.800000 0.600000 ;
    END
  END pmem_out2[56]
  PIN pmem_out2[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.200000 0.000000 405.400000 0.600000 ;
    END
  END pmem_out2[55]
  PIN pmem_out2[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.800000 0.000000 405.000000 0.600000 ;
    END
  END pmem_out2[54]
  PIN pmem_out2[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.400000 0.000000 404.600000 0.600000 ;
    END
  END pmem_out2[53]
  PIN pmem_out2[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.000000 0.000000 404.200000 0.600000 ;
    END
  END pmem_out2[52]
  PIN pmem_out2[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.600000 0.000000 403.800000 0.600000 ;
    END
  END pmem_out2[51]
  PIN pmem_out2[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.200000 0.000000 403.400000 0.600000 ;
    END
  END pmem_out2[50]
  PIN pmem_out2[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.800000 0.000000 403.000000 0.600000 ;
    END
  END pmem_out2[49]
  PIN pmem_out2[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.400000 0.000000 402.600000 0.600000 ;
    END
  END pmem_out2[48]
  PIN pmem_out2[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.000000 0.000000 402.200000 0.600000 ;
    END
  END pmem_out2[47]
  PIN pmem_out2[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.600000 0.000000 401.800000 0.600000 ;
    END
  END pmem_out2[46]
  PIN pmem_out2[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.200000 0.000000 401.400000 0.600000 ;
    END
  END pmem_out2[45]
  PIN pmem_out2[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.800000 0.000000 401.000000 0.600000 ;
    END
  END pmem_out2[44]
  PIN pmem_out2[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.400000 0.000000 400.600000 0.600000 ;
    END
  END pmem_out2[43]
  PIN pmem_out2[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.000000 0.000000 400.200000 0.600000 ;
    END
  END pmem_out2[42]
  PIN pmem_out2[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.600000 0.000000 399.800000 0.600000 ;
    END
  END pmem_out2[41]
  PIN pmem_out2[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.200000 0.000000 399.400000 0.600000 ;
    END
  END pmem_out2[40]
  PIN pmem_out2[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.800000 0.000000 399.000000 0.600000 ;
    END
  END pmem_out2[39]
  PIN pmem_out2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.400000 0.000000 398.600000 0.600000 ;
    END
  END pmem_out2[38]
  PIN pmem_out2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.000000 0.000000 398.200000 0.600000 ;
    END
  END pmem_out2[37]
  PIN pmem_out2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.600000 0.000000 397.800000 0.600000 ;
    END
  END pmem_out2[36]
  PIN pmem_out2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.200000 0.000000 397.400000 0.600000 ;
    END
  END pmem_out2[35]
  PIN pmem_out2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.800000 0.000000 397.000000 0.600000 ;
    END
  END pmem_out2[34]
  PIN pmem_out2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.400000 0.000000 396.600000 0.600000 ;
    END
  END pmem_out2[33]
  PIN pmem_out2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.000000 0.000000 396.200000 0.600000 ;
    END
  END pmem_out2[32]
  PIN pmem_out2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.600000 0.000000 395.800000 0.600000 ;
    END
  END pmem_out2[31]
  PIN pmem_out2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.200000 0.000000 395.400000 0.600000 ;
    END
  END pmem_out2[30]
  PIN pmem_out2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.800000 0.000000 395.000000 0.600000 ;
    END
  END pmem_out2[29]
  PIN pmem_out2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.400000 0.000000 394.600000 0.600000 ;
    END
  END pmem_out2[28]
  PIN pmem_out2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.000000 0.000000 394.200000 0.600000 ;
    END
  END pmem_out2[27]
  PIN pmem_out2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.600000 0.000000 393.800000 0.600000 ;
    END
  END pmem_out2[26]
  PIN pmem_out2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.200000 0.000000 393.400000 0.600000 ;
    END
  END pmem_out2[25]
  PIN pmem_out2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.800000 0.000000 393.000000 0.600000 ;
    END
  END pmem_out2[24]
  PIN pmem_out2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.400000 0.000000 392.600000 0.600000 ;
    END
  END pmem_out2[23]
  PIN pmem_out2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.000000 0.000000 392.200000 0.600000 ;
    END
  END pmem_out2[22]
  PIN pmem_out2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.600000 0.000000 391.800000 0.600000 ;
    END
  END pmem_out2[21]
  PIN pmem_out2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.200000 0.000000 391.400000 0.600000 ;
    END
  END pmem_out2[20]
  PIN pmem_out2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.800000 0.000000 391.000000 0.600000 ;
    END
  END pmem_out2[19]
  PIN pmem_out2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.400000 0.000000 390.600000 0.600000 ;
    END
  END pmem_out2[18]
  PIN pmem_out2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.000000 0.000000 390.200000 0.600000 ;
    END
  END pmem_out2[17]
  PIN pmem_out2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.600000 0.000000 389.800000 0.600000 ;
    END
  END pmem_out2[16]
  PIN pmem_out2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.200000 0.000000 389.400000 0.600000 ;
    END
  END pmem_out2[15]
  PIN pmem_out2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.800000 0.000000 389.000000 0.600000 ;
    END
  END pmem_out2[14]
  PIN pmem_out2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.400000 0.000000 388.600000 0.600000 ;
    END
  END pmem_out2[13]
  PIN pmem_out2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.000000 0.000000 388.200000 0.600000 ;
    END
  END pmem_out2[12]
  PIN pmem_out2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.600000 0.000000 387.800000 0.600000 ;
    END
  END pmem_out2[11]
  PIN pmem_out2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.200000 0.000000 387.400000 0.600000 ;
    END
  END pmem_out2[10]
  PIN pmem_out2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.800000 0.000000 387.000000 0.600000 ;
    END
  END pmem_out2[9]
  PIN pmem_out2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.400000 0.000000 386.600000 0.600000 ;
    END
  END pmem_out2[8]
  PIN pmem_out2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.000000 0.000000 386.200000 0.600000 ;
    END
  END pmem_out2[7]
  PIN pmem_out2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.600000 0.000000 385.800000 0.600000 ;
    END
  END pmem_out2[6]
  PIN pmem_out2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.200000 0.000000 385.400000 0.600000 ;
    END
  END pmem_out2[5]
  PIN pmem_out2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.800000 0.000000 385.000000 0.600000 ;
    END
  END pmem_out2[4]
  PIN pmem_out2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.400000 0.000000 384.600000 0.600000 ;
    END
  END pmem_out2[3]
  PIN pmem_out2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.000000 0.000000 384.200000 0.600000 ;
    END
  END pmem_out2[2]
  PIN pmem_out2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.600000 0.000000 383.800000 0.600000 ;
    END
  END pmem_out2[1]
  PIN pmem_out2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.200000 0.000000 383.400000 0.600000 ;
    END
  END pmem_out2[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 766.400000 765.200000 ;
    LAYER M2 ;
      RECT 0.000000 0.700000 766.400000 765.200000 ;
      RECT 459.900000 0.000000 766.400000 0.700000 ;
      RECT 0.000000 0.000000 306.300000 0.700000 ;
    LAYER M3 ;
      RECT 0.000000 407.600000 766.400000 765.200000 ;
      RECT 0.700000 357.200000 766.400000 407.600000 ;
      RECT 0.000000 0.000000 766.400000 357.200000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 766.400000 765.200000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 766.400000 765.200000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 766.400000 765.200000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 766.400000 765.200000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 766.400000 765.200000 ;
  END
END fullchip

END LIBRARY
